module siguelineas ( 
	si,
	sd,
	mi,
	md
	) ;

input  si;
input  sd;
inout  mi;
inout  md;

module tubo1 ( 
	clk,
	reset,
	q
	) ;

input  clk;
input  reset;
inout [6:0] q;

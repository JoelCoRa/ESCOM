module mario ( 
	clk,
	sw,
	q
	) ;

input  clk;
input  sw;
inout [2:0] q;

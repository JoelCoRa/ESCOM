module piso ( 
	clk,
	q
	) ;

input  clk;
inout  q;

module escenario ( 
	clk,
	output,
	reset
	) ;

input  clk;
inout [6:0] output;
input  reset;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DSD IS
PORT(
    D0,D1,D2,D3,D4,D5,D6,D7,D8,D9:IN STD_LOGIC;
	SAL0,SAL1,SAL2,SAL3,SAL4,SAL5,SAL6,SAL7,SAL8,SAL9: OUT STD_LOGIC);

ATTRIBUTE PIN_NUMBERS OF DSD: ENTITY IS
"D0:1 D1:2 D2:3 D3:4 D4:5 D5:6 D6:7 D7:8 D8:9 SAL0:23 SAL1:22 SAL2:21 SAL3:20 SAL4:19 SAL5:18 SAL6:17 SAL7:16 SAL8:15";
END ENTITY;
ARCHITECTURE ENCIENDE OF DSD IS
BEGIN
  SAL0<=D0;
  SAL1<=D1;
  SAL2<=D2;
  SAL3<=D3;
  SAL4<=D4;
  SAL5<=D5;
  SAL6<=D6;
  SAL7<=D7;
  SAL8<=D8;
  SAL9<=D9;
END ENCIENDE;

